-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.0 Build 184 04/29/2009 Service Pack 1 SJ Web Edition
-- Created on Mon May 17 19:52:14 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FIFOcontrol IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        rdempty_1 : IN STD_LOGIC := '0';
        wrfull_1 : IN STD_LOGIC := '0';
        wrfull_2 : IN STD_LOGIC := '0';
        wr1 : OUT STD_LOGIC;
        wr2 : OUT STD_LOGIC;
        rd1 : OUT STD_LOGIC;
        rd2 : OUT STD_LOGIC
    );
END FIFOcontrol;

ARCHITECTURE BEHAVIOR OF FIFOcontrol IS
    TYPE type_fstate IS (initial_1,w1,r1w2,w1r2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= initial_1;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,rdempty_1,wrfull_1,wrfull_2)
    BEGIN
        wr1 <= '0';
        wr2 <= '0';
        rd1 <= '0';
        rd2 <= '0';
        CASE fstate IS
            WHEN initial_1 =>
                IF ((rdempty_1 = '1')) THEN
                    reg_fstate <= w1;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= initial_1;
                END IF;

                wr2 <= '0';

                rd2 <= '0';

                wr1 <= '1';

                rd1 <= '0';
            WHEN w1 =>
                IF ((wrfull_1 = '1')) THEN
                    reg_fstate <= r1w2;
                ELSE
                    reg_fstate <= w1;
                END IF;

                wr2 <= '0';

                rd2 <= '0';

                wr1 <= '1';

                rd1 <= '0';
            WHEN r1w2 =>
                IF ((wrfull_2 = '1')) THEN
                    reg_fstate <= w1r2;
                ELSE
                    reg_fstate <= r1w2;
                END IF;

                wr2 <= '1';

                rd2 <= '0';

                wr1 <= '0';

                rd1 <= '1';
            WHEN w1r2 =>
                IF ((wrfull_1 = '1')) THEN
                    reg_fstate <= r1w2;
                ELSE
                    reg_fstate <= w1r2;
                END IF;

                wr2 <= '0';

                rd2 <= '1';

                wr1 <= '1';

                rd1 <= '0';
            WHEN OTHERS => 
                wr1 <= 'X';
                wr2 <= 'X';
                rd1 <= 'X';
                rd2 <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
